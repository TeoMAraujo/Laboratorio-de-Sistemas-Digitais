library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity arithmetic_control is
    port (
        OPCODE   : in    std_logic_vector(2 downto 0);
        OPERAND1 : in    std_logic_vector(7 downto 0);
        OPERAND2 : in    std_logic_vector(2 downto 0);
        CLK      : in    std_logic;
        RST      : in    std_logic; 
        OUTP     : out   std_logic_vector(7 downto 0);
        ADDR     : out   std_logic_vector(2 downto 0);
        DATA     : inout std_logic_vector(7 downto 0);
        READW    : out   std_logic
    );
end arithmetic_control;

architecture structural of arithmetic_control is
    signal toALUB              : std_logic_vector(7 downto 0) := (others => '0');
    signal toMuxA              : std_logic_vector(2 downto 0) := (others => '0');
    signal toMuxB              : std_logic_vector(7 downto 0);
    alias toMuxBAddr is toMuxB (2 downto 0);
    
    signal toMuxS              : std_logic := '0';
    signal toDemuxA            : std_logic_vector(7 downto 0) := (others => '0');
    signal toDemuxSel_read_dff : std_logic := '0';
    signal toALUS_Comparator   : std_logic_vector(2 downto 0) := (others => '0');
    signal demux_to_data_bus   : std_logic_vector(7 downto 0);
    signal opcode_pipe1        : std_logic_vector(2 downto 0) := (others => '0');
    
    signal demux_select_inv    : std_logic; 

begin
    -- CYCLE 1 
    U_DFF1: entity work.D_flip_flop
        generic map (W => 3) -- NOTE: Removed incorrect semicolon here
        port map (D => OPCODE, CLK => CLK, RST => RST, Q => toALUS_Comparator, Qn => open);

    U_DFF2: entity work.D_flip_flop
        generic map (W => 8)
        port map (D => OPERAND1, CLK => CLK, RST => RST, Q => toDemuxA, Qn => open);

    U_DFF3: entity work.D_flip_flop
        generic map (W => 3)
        port map (D => OPERAND2, CLK => CLK, RST => RST, Q => toMuxA, Qn => open);

    U_COMP: entity work.comparator
        generic map (W => 3)
        port map (A => toALUS_Comparator, B => "000", equal => toDemuxSel_Read_dff);

    demux_select_inv <= not toDemuxSel_Read_dff;

    U_DEMUX: entity work.Demux_1x2
        generic map (W => 8)
        port map (
            A  => toDemuxA, 
            S  => demux_select_inv, 
            Y0 => demux_to_data_bus, 
            Y1 => toMuxB
        );

    DATA <= demux_to_data_bus when toDemuxSel_Read_dff = '1' else (others => 'Z');
    
    toMuxS <= toDemuxSel_Read_dff; 

    U_MUX: entity work.Mux_2x1
        generic map(W => 3)
        port map (A => toMuxBAddr, B => toMuxA, S => toMuxS, Y => ADDR);

    -- CYCLE 2
    U_DFF5: entity work.D_flip_flop
        generic map (W => 8)
        port map (D => DATA, CLK => CLK, RST => RST, Q => toALUB, Qn => open);

    U_DFFALU1: entity work.D_flip_flop
        generic map (W => 3)
        port map (D => toALUS_Comparator, CLK => CLK, RST => RST, Q => opcode_pipe1, Qn => open);

    U_ALU: entity work.ALU
        generic map (W => 8)
        port map (
            A      => DATA,            
            B      => toALUB,         
            opcode => opcode_pipe1, 
            Y      => OUTP
        );
        
    READW <= toDemuxSel_Read_dff;
end structural;
